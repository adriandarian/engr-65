** Profile: "SCHEMATIC1-lab6"  [ C:\Users\adarian\Documents\ucmerced-coursework\engr-65\Labs\Lab-6\Lab6-PSpiceFiles\SCHEMATIC1\lab6.sim ] 

** Creating circuit file "lab6.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
* From [PSPICE NETLIST] section of C:\SPB_DATA\cdssetup\OrCAD_PSpice\17.4.0\PSpice.ini file:
.lib "nom.lib" 

*Analysis directives: 
.TRAN  0 40ms 0 5us 
.OPTIONS ADVCONV
.PROBE64 N([N14434])
.PROBE64 N([N14438])
.INC "..\SCHEMATIC1.net" 


.END
